/*
*  File            :   nf_csr.svh
*  Autor           :   Vlasov D.V.
*  Data            :   2019.05.16
*  Language        :   SystemVerilog
*  Description     :   This is CSR constants
*  Copyright(c)    :   2018 - 2019 Vlasov D.V.
*/

`define USTATUS_A   12'h000
`define UIE_A       12'h004
`define UTVEC_A     12'h005  
`define MCYCLE_A    12'hB00
