/*
*  File            :   nf_hazard_unit.sv
*  Autor           :   Vlasov D.V.
*  Data            :   2019.01.10
*  Language        :   SystemVerilog
*  Description     :   This is hazard unit constants
*  Copyright(c)    :   2018 - 2019 Vlasov D.V.
*/

`define     HU_BP_NONE  2'b00
`define     HU_BP_MEM   2'b01
`define     HU_BP_WB    2'b10
