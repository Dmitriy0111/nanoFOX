/*
*  File            :   nf_tb.svh
*  Autor           :   Vlasov D.V.
*  Data            :   2018.11.28
*  Language        :   SystemVerilog
*  Description     :   This is testbench header for cpu unit
*  Copyright(c)    :   2018 - 2019 Vlasov D.V.
*/

// enable debug instruction messages
`define debug_lev0  1
// enable logging
`define log_en      1
// enable logging
`define log_html    1
