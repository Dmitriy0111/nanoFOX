/*
*  File            :   nf_tb.svh
*  Autor           :   Vlasov D.V.
*  Data            :   2018.11.28
*  Language        :   SystemVerilog
*  Description     :   This is testbench header for cpu unit
*  Copyright(c)    :   2018 Vlasov D.V.
*/

`define debug_lev0
